* AD8217 SPICE Macro-model
* Description: Zero-Drift Current Shunt Monitor
* Generic Desc: 4.5V to 80V operation, high side current sensing
* Developed by: DK
* Revision History:
* 1.0 (9/2012) - DK - initial release
* 1.1 (10/2012) - DK - netlist change
* Copyright 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html
* for License Statement. Use of this model indicates your acceptance
* of the terms and provisions in the License Statement.
*
*
* Not Modeled:
* Temperature effects
* PSRR vs Frequency
*
* Parameters modeled include:
* CMRR vs Frequency
* VOS (RTI)
* Bandwidth
* Gain Error
* Voltage Spectral Noise: 110nV/rt hz at 1kHz
* Output Impedance: 2 ohms
* Common Mode Range: 4.5V to 80V
*
* END Notes
* Maximum output voltage limited to 5.6V
*
* Node Assignments
*                 noninverting input
*                 |   inverting input
*                 |   |   ground
*                 |   |   |   output
*                 |   |   |   |
.SUBCKT AD8217  +IN -IN GND OUT

*** Input Stage ***
Q1 3 1 7. 0 NPN
Q2 4 2 8 0 NPN
R1 +IN 3 1129
R2 +IN 4 1129
R3 7. 9 1e3
R4 8 9 1e3
I1 9 GND 400E-6
Ibp +IN GND 157E-6
Ibn -IN GND 16E-6

*** Input and Feedback Resistors ***
EOS 5 1 poly(1) (201,GND) 0 -1
R9 5 +IN 75e3
R10 GND 5 1.5e6
R11 -IN 2 75.045e3
R12 20 2 1.5e6

*** 1st Stage ***
D1 100 6 DZENER2
G1 100 10 1 2 .001
D2 10 6 DZENER1
R8 10 100 200e3

*** 2nd Stage ***
G2 100 20 10 100 .005
R7 20 100 1E6
C1 20 100 11.68E-9

*** Internal Reference ***
E1 100 0 7 0 1
R5 +IN 7 100e3
R6 7 GND 100e3

**** zero-pole stage
*G4 100 30 20 100 .59e-6
G4 100 30 20 100 .588e-6
R14 30 35 1e6
R16 35 100 1.7e6
L1 30 35 .65

**** 1st pole stage
G3 100 40 30 100 1e-6
R13 40 100 1E6
C2 40 100 186e-15

**** 2nd pole stage
G5 100 45 40 100 1e-6
R15 45 100 1E6
C3 45 100 186e-15


*** Spectral Noise ***
VN GND 190 .65
DN 190 200 DNOISE
RN 200 GND 1
VM GND 200 0
FN GND 201 VM 1
RZ 201 GND 1

*** CMRR ***
GCMR 500 0 505 0 .3e-9
RCM1 500 501 549e6
LCMR 500 501 80
RCM2 501 0 1e6

GCM2 600 0 500 0 .85e-6
RCM3 600 0 1e6
CCM2 600 0 655e-15

RCMR1 +IN 505 10e6
RCMR2 505 -IN 10e6

*** Clamp
D3 11 20 D
V7 11 0 0

*** Output Stage ***
EAVG AVG GND Value={ ((V(+IN) + V(-IN))*0.5 )}
E01 60 0 Value={ IF( V(45) > 5.6, 5.6 , IF( V(45) < 5.6, V(45) - .002, V(45) )) }
E02 65 0 Value={ IF( V(AVG) > 80, 5.6 , IF( V(AVG) < 4.5, 0, V(60) )) }
EO3 70 0 value = { (V(65) + V(600)) }

*** Output Resistance
Rout 70 OUT 2

*** Output Current limiting
Et 71 0 70 OUT 20
Qc 45 71 72 0 NPN
Rb 72 0 10

.model D D(IS=5.950e-006 N=4.031e+000 RS=2.677e-002)
.model DZENER1 D(BV=2V, IS=1E-14, IBV=1E-3)
.model DZENER2 D(BV=2V, IS=1E-14, IBV=1E-3)
.model DNOISE D(AF=0, KF=0.0195e-10.5)
.model DILIM D(IS=1E-15)
.model NPN NPN

.ends